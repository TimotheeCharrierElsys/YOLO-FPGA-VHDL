library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

library LIB_RTL;
use LIB_RTL.types_pkg.all;

entity conv_tb is
end;

architecture conv_tb_arch of conv_tb is
    -- Clock period
    constant i_clk_period : time := 5 ns;
    -- Generics
    constant BITWIDTH       : integer := 8;
    constant INPUT_SIZE     : integer := 64;
    constant CHANNEL_NUMBER : integer := 3;
    constant KERNEL_SIZE    : integer := 3;
    constant KERNEL_NUMBER  : integer := 3;
    constant PADDING        : integer := 1;
    constant STRIDE         : integer := 1;
    -- Ports
    signal clock        : std_logic                                                                                                                                           := '0';
    signal reset_n      : std_logic                                                                                                                                           := '0';
    signal i_sys_enable : std_logic                                                                                                                                           := '0';
    signal i_data_valid : std_logic                                                                                                                                           := '0';
    signal i_data       : t_volume(CHANNEL_NUMBER - 1 downto 0)(INPUT_SIZE - 1 downto 0)(INPUT_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0)                                      := (others => (others => (others => (others => '0'))));
    signal i_kernel     : t_input_feature(KERNEL_NUMBER - 1 downto 0)(CHANNEL_NUMBER - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0) := (others => (others => (others => (others => (others => '0')))));
    signal i_bias       : t_vec(KERNEL_NUMBER - 1 downto 0)(BITWIDTH - 1 downto 0);
    signal o_data       : t_volume(KERNEL_NUMBER - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)(2 * BITWIDTH - 1 downto 0);
    signal o_data_valid : std_logic;

    -- File variables
    file output_file : text;

    component conv
        generic (
            BITWIDTH       : integer;
            INPUT_SIZE     : integer;
            CHANNEL_NUMBER : integer;
            KERNEL_SIZE    : integer;
            KERNEL_NUMBER  : integer;
            PADDING        : integer;
            STRIDE         : integer
        );
        port (
            clock        : in std_logic;
            reset_n      : in std_logic;
            i_sys_enable : in std_logic;
            i_data_valid : in std_logic;
            i_data       : in t_volume(CHANNEL_NUMBER - 1 downto 0)(INPUT_SIZE - 1 downto 0)(INPUT_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0);
            i_kernel     : in t_input_feature(KERNEL_NUMBER - 1 downto 0)(CHANNEL_NUMBER - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0);
            i_bias       : in t_vec(KERNEL_NUMBER - 1 downto 0)(BITWIDTH - 1 downto 0);
            o_data       : out t_volume(KERNEL_NUMBER - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)(2 * BITWIDTH - 1 downto 0);
            o_data_valid : out std_logic
        );
    end component;

begin

    UUT : conv
    generic map(
        BITWIDTH       => BITWIDTH,
        INPUT_SIZE     => INPUT_SIZE,
        CHANNEL_NUMBER => CHANNEL_NUMBER,
        KERNEL_SIZE    => KERNEL_SIZE,
        KERNEL_NUMBER  => KERNEL_NUMBER,
        PADDING        => PADDING,
        STRIDE         => STRIDE
    )
    port map(
        clock        => clock,
        reset_n      => reset_n,
        i_sys_enable => i_sys_enable,
        i_data_valid => i_data_valid,
        i_data       => i_data,
        i_kernel     => i_kernel,
        i_bias       => i_bias,
        o_data       => o_data,
        o_data_valid => o_data_valid
    );

    i_bias <= (others => std_logic_vector(to_signed(0, BITWIDTH)));

    -- Clock generation
    clock <= not clock after i_clk_period / 2;

    -------------------------------------------------------------------------------------
    -- TEST PROCESS
    -------------------------------------------------------------------------------------
    stimulus : process
        variable line_buffer : line;
    begin
        -- Reset the system
        reset_n      <= '0';
        i_data_valid <= '0';
        wait for i_clk_period;
        reset_n      <= '1';
        i_sys_enable <= '1';

        i_data(0) <= (
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(108, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(129, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(139, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(165, 8))),
        (std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(194, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(172, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(159, 8))),
        (std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(185, 8))),
        (std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(183, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(181, 8))),
        (std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(161, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(255, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(105, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(249, 8)), std_logic_vector(to_signed(249, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(41, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(244, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(241, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(237, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8))),
        (std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(238, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8))),
        (std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(238, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(235, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8))),
        (std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8))),
        (std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(25, 8))),
        (std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(15, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8))),
        (std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(40, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(237, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(38, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(235, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(79, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(244, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(235, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(242, 8)), std_logic_vector(to_signed(235, 8)), std_logic_vector(to_signed(201, 8))),
        (std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(238, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(225, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(237, 8)), std_logic_vector(to_signed(250, 8)), std_logic_vector(to_signed(231, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(243, 8)), std_logic_vector(to_signed(238, 8))),
        (std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(241, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(238, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(240, 8))),
        (std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(228, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(253, 8)), std_logic_vector(to_signed(255, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(241, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(237, 8))),
        (std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(242, 8)), std_logic_vector(to_signed(252, 8)), std_logic_vector(to_signed(245, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(235, 8)), std_logic_vector(to_signed(245, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(235, 8)), std_logic_vector(to_signed(248, 8)), std_logic_vector(to_signed(232, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(230, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(203, 8))),
        (std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(237, 8)), std_logic_vector(to_signed(236, 8)), std_logic_vector(to_signed(237, 8)), std_logic_vector(to_signed(235, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(249, 8)), std_logic_vector(to_signed(240, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(234, 8)), std_logic_vector(to_signed(238, 8)), std_logic_vector(to_signed(233, 8)), std_logic_vector(to_signed(229, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(189, 8))),
        (std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(221, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(226, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(242, 8)), std_logic_vector(to_signed(250, 8)), std_logic_vector(to_signed(239, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(148, 8))),
        (std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(158, 8))),
        (std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(162, 8))),
        (std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(174, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(221, 8))),
        (std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(222, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(201, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(218, 8)), std_logic_vector(to_signed(225, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(186, 8))),
        (std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(212, 8)), std_logic_vector(to_signed(211, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(223, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(214, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(227, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(224, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(54, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(217, 8)), std_logic_vector(to_signed(213, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8))),
        (std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(6, 8))),
        (std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(43, 8))),
        (std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(40, 8))),
        (std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(39, 8))),
        (std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8))),
        (std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8))),
        (std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(37, 8))),
        (std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(32, 8))),
        (std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(32, 8))),
        (std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(29, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(46, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(30, 8))),
        (std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(26, 8))),
        (std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(17, 8))),
        (std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8))),
        (std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(17, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(21, 8)))
        );
        i_data(1) <= (
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(62, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(86, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(115, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(136, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(102, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(65, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(80, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(77, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(92, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(103, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(219, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(73, 8))),
        (std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(208, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(209, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(30, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(41, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(30, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(207, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(206, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8))),
        (std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8))),
        (std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(34, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(20, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8))),
        (std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8))),
        (std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(203, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(19, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(195, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(50, 8))),
        (std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(204, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(161, 8))),
        (std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(172, 8))),
        (std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(176, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(179, 8))),
        (std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(180, 8))),
        (std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(198, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(155, 8))),
        (std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(152, 8))),
        (std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(197, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(122, 8))),
        (std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(132, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(128, 8))),
        (std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(126, 8))),
        (std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(159, 8))),
        (std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(136, 8))),
        (std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(133, 8))),
        (std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(19, 8))),
        (std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(36, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(6, 8))),
        (std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(36, 8))),
        (std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(30, 8))),
        (std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(29, 8))),
        (std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(33, 8))),
        (std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(33, 8))),
        (std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(27, 8))),
        (std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(24, 8))),
        (std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(24, 8))),
        (std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(22, 8))),
        (std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(42, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(27, 8))),
        (std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(26, 8))),
        (std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(18, 8))),
        (std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8))),
        (std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(19, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(23, 8)))
        );
        i_data(2) <= (
        (std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(35, 8))),
        (std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(53, 8))),
        (std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(54, 8))),
        (std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(66, 8))),
        (std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(72, 8))),
        (std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(32, 8))),
        (std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(1, 8))),
        (std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(23, 8))),
        (std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(35, 8))),
        (std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(62, 8))),
        (std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(81, 8))),
        (std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(58, 8))),
        (std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(21, 8))),
        (std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(25, 8))),
        (std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8))),
        (std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(196, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(28, 8))),
        (std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(210, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(30, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(220, 8)), std_logic_vector(to_signed(216, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8))),
        (std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(215, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(22, 8))),
        (std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(22, 8))),
        (std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(20, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(73, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(22, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8))),
        (std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(199, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8))),
        (std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(68, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(16, 8))),
        (std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(30, 8))),
        (std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(200, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8))),
        (std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(201, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(5, 8))),
        (std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(205, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(32, 8))),
        (std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(202, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(135, 8))),
        (std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(132, 8))),
        (std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(191, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(137, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(166, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(151, 8))),
        (std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(161, 8))),
        (std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(141, 8))),
        (std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(187, 8)), std_logic_vector(to_signed(190, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(134, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(185, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(148, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(95, 8))),
        (std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(97, 8))),
        (std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(140, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(82, 8))),
        (std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(181, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(77, 8))),
        (std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(180, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(183, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(112, 8))),
        (std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(188, 8)), std_logic_vector(to_signed(194, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(157, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(96, 8))),
        (std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(189, 8)), std_logic_vector(to_signed(174, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(158, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(102, 8))),
        (std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(179, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(193, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(172, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(0, 8))),
        (std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(66, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(192, 8)), std_logic_vector(to_signed(178, 8)), std_logic_vector(to_signed(184, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(161, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(19, 8))),
        (std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(182, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(186, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(165, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(142, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(0, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(70, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(177, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(159, 8)), std_logic_vector(to_signed(155, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(26, 8))),
        (std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(62, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(170, 8)), std_logic_vector(to_signed(175, 8)), std_logic_vector(to_signed(164, 8)), std_logic_vector(to_signed(171, 8)), std_logic_vector(to_signed(163, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(133, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(122, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(119, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(137, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(21, 8))),
        (std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(162, 8)), std_logic_vector(to_signed(176, 8)), std_logic_vector(to_signed(169, 8)), std_logic_vector(to_signed(160, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(153, 8)), std_logic_vector(to_signed(147, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(136, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(20, 8))),
        (std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(59, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(60, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(168, 8)), std_logic_vector(to_signed(151, 8)), std_logic_vector(to_signed(156, 8)), std_logic_vector(to_signed(152, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(128, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(111, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(24, 8))),
        (std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(173, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(154, 8)), std_logic_vector(to_signed(150, 8)), std_logic_vector(to_signed(146, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(125, 8)), std_logic_vector(to_signed(120, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(103, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(23, 8))),
        (std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(63, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(130, 8)), std_logic_vector(to_signed(167, 8)), std_logic_vector(to_signed(149, 8)), std_logic_vector(to_signed(144, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(134, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(123, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(71, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(17, 8))),
        (std_logic_vector(to_signed(64, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(65, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(145, 8)), std_logic_vector(to_signed(141, 8)), std_logic_vector(to_signed(139, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(131, 8)), std_logic_vector(to_signed(126, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(112, 8)), std_logic_vector(to_signed(104, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(13, 8))),
        (std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(82, 8)), std_logic_vector(to_signed(46, 8)), std_logic_vector(to_signed(53, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(143, 8)), std_logic_vector(to_signed(138, 8)), std_logic_vector(to_signed(135, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(124, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(110, 8)), std_logic_vector(to_signed(102, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(13, 8))),
        (std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(107, 8)), std_logic_vector(to_signed(113, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(132, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(118, 8)), std_logic_vector(to_signed(116, 8)), std_logic_vector(to_signed(105, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(100, 8)), std_logic_vector(to_signed(97, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(94, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(5, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(12, 8))),
        (std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(61, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(84, 8)), std_logic_vector(to_signed(127, 8)), std_logic_vector(to_signed(129, 8)), std_logic_vector(to_signed(117, 8)), std_logic_vector(to_signed(115, 8)), std_logic_vector(to_signed(114, 8)), std_logic_vector(to_signed(108, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(69, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(31, 8))),
        (std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(121, 8)), std_logic_vector(to_signed(106, 8)), std_logic_vector(to_signed(89, 8)), std_logic_vector(to_signed(101, 8)), std_logic_vector(to_signed(98, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(95, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(90, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(91, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(93, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(87, 8)), std_logic_vector(to_signed(96, 8)), std_logic_vector(to_signed(72, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(18, 8))),
        (std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(109, 8)), std_logic_vector(to_signed(99, 8)), std_logic_vector(to_signed(92, 8)), std_logic_vector(to_signed(88, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(79, 8)), std_logic_vector(to_signed(81, 8)), std_logic_vector(to_signed(74, 8)), std_logic_vector(to_signed(83, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(16, 8))),
        (std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(40, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(52, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(6, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(86, 8)), std_logic_vector(to_signed(85, 8)), std_logic_vector(to_signed(80, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(77, 8)), std_logic_vector(to_signed(75, 8)), std_logic_vector(to_signed(76, 8)), std_logic_vector(to_signed(78, 8)), std_logic_vector(to_signed(67, 8)), std_logic_vector(to_signed(54, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(1, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(3, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(4, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(10, 8))),
        (std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(31, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(36, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(58, 8)), std_logic_vector(to_signed(55, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(33, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(28, 8))),
        (std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(51, 8)), std_logic_vector(to_signed(47, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(37, 8)), std_logic_vector(to_signed(44, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(17, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(16, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(0, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(14, 8))),
        (std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(48, 8)), std_logic_vector(to_signed(57, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(56, 8)), std_logic_vector(to_signed(50, 8)), std_logic_vector(to_signed(49, 8)), std_logic_vector(to_signed(41, 8)), std_logic_vector(to_signed(18, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(43, 8)), std_logic_vector(to_signed(38, 8)), std_logic_vector(to_signed(45, 8)), std_logic_vector(to_signed(42, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(22, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(27, 8)), std_logic_vector(to_signed(21, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(11, 8)), std_logic_vector(to_signed(7, 8)), std_logic_vector(to_signed(9, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(25, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(32, 8)), std_logic_vector(to_signed(23, 8)), std_logic_vector(to_signed(34, 8)), std_logic_vector(to_signed(39, 8)), std_logic_vector(to_signed(20, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(30, 8)), std_logic_vector(to_signed(29, 8)), std_logic_vector(to_signed(2, 8)), std_logic_vector(to_signed(26, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(13, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(8, 8)), std_logic_vector(to_signed(10, 8)), std_logic_vector(to_signed(14, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(28, 8)), std_logic_vector(to_signed(15, 8)), std_logic_vector(to_signed(35, 8)), std_logic_vector(to_signed(12, 8)), std_logic_vector(to_signed(19, 8)), std_logic_vector(to_signed(24, 8)), std_logic_vector(to_signed(18, 8)))
        );

        i_kernel(0)(0) <= (others => (others => std_logic_vector(to_signed(1, BITWIDTH))));
        i_kernel(0)(1) <= (others => (others => std_logic_vector(to_signed(1, BITWIDTH))));
        i_kernel(0)(2) <= (others => (others => std_logic_vector(to_signed(1, BITWIDTH))));

        i_kernel(1)(0) <= ((std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH))));
        i_kernel(1)(1) <= ((std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH))));
        i_kernel(1)(2) <= ((std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH))));
        
        i_kernel(2)(0) <= ((std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH))));
        i_kernel(2)(1) <= ((std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH))));
        i_kernel(2)(2) <= ((std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH))),
        (std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(0, BITWIDTH)), std_logic_vector(to_signed(1, BITWIDTH))));

        wait for i_clk_period/2;
        i_data_valid <= '1';
        wait for i_clk_period;
        i_data_valid <= '0';

        -- Open the file
        file_open(output_file, "conv_output_results.txt", write_mode);

        -- Wait for output to be valid and write to file
        wait until o_data_valid = '1';
        for k in 0 to KERNEL_NUMBER - 1 loop
            for i in 0 to ((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1) loop
                for j in 0 to ((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1) loop
                    write(line_buffer, o_data(k)(i)(j));
                    writeline(output_file, line_buffer);
                end loop;
            end loop;
        end loop;

        -- Close the file
        file_close(output_file);

        -- End simulation
        wait;

    end process stimulus;
end conv_tb_arch;

configuration conv_tb_conf of conv_tb is
    for conv_tb_arch
        for UUT : conv
            use configuration LIB_RTL.conv_fc_conf;
        end for;
    end for;
end configuration conv_tb_conf;