library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

library LIB_RTL;
use LIB_RTL.types_pkg.all;

entity conv2d_tb is
end;

architecture conv2d_tb_arch of conv2d_tb is
    -- Clock period
    constant i_clk_period : time := 5 ns;
    -- Generics
    constant BITWIDTH       : integer := 16;
    constant INPUT_SIZE     : integer := 64;
    constant CHANNEL_NUMBER : integer := 3;
    constant KERNEL_SIZE    : integer := 3;
    constant KERNEL_NUMBER  : integer := 13;
    constant PADDING        : integer := 1;
    constant STRIDE         : integer := 1;
    -- Ports
    signal clock        : std_logic                                                                                                                                           := '0';
    signal reset_n      : std_logic                                                                                                                                           := '0';
    signal i_sys_enable : std_logic                                                                                                                                           := '0';
    signal i_data_valid : std_logic                                                                                                                                           := '0';
    signal i_data       : t_volume(CHANNEL_NUMBER - 1 downto 0)(INPUT_SIZE - 1 downto 0)(INPUT_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0)                                      := (others => (others => (others => (others => '0'))));
    signal i_kernel     : t_input_feature(KERNEL_NUMBER - 1 downto 0)(CHANNEL_NUMBER - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0) := (others => (others => (others => (others => (others => '0')))));
    signal i_bias       : t_vec(KERNEL_NUMBER - 1 downto 0)(BITWIDTH - 1 downto 0);
    signal o_data       : t_volume(KERNEL_NUMBER - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)(2 * BITWIDTH - 1 downto 0);
    signal o_data_valid : std_logic;

    -- File variables
    file output_file : text;

    component conv2d
        generic (
            BITWIDTH       : integer;
            INPUT_SIZE     : integer;
            CHANNEL_NUMBER : integer;
            KERNEL_SIZE    : integer;
            KERNEL_NUMBER  : integer;
            PADDING        : integer;
            STRIDE         : integer
        );
        port (
            clock        : in std_logic;
            reset_n      : in std_logic;
            i_sys_enable : in std_logic;
            i_data_valid : in std_logic;
            i_data       : in t_volume(CHANNEL_NUMBER - 1 downto 0)(INPUT_SIZE - 1 downto 0)(INPUT_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0);
            i_kernel     : in t_input_feature(KERNEL_NUMBER - 1 downto 0)(CHANNEL_NUMBER - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(KERNEL_SIZE - 1 downto 0)(BITWIDTH - 1 downto 0);
            i_bias       : in t_vec(KERNEL_NUMBER - 1 downto 0)(BITWIDTH - 1 downto 0);
            o_data       : out t_volume(KERNEL_NUMBER - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1 downto 0)(2 * BITWIDTH - 1 downto 0);
            o_data_valid : out std_logic
        );
    end component;

begin

    UUT : conv2d
    generic map(
        BITWIDTH       => BITWIDTH,
        INPUT_SIZE     => INPUT_SIZE,
        CHANNEL_NUMBER => CHANNEL_NUMBER,
        KERNEL_SIZE    => KERNEL_SIZE,
        KERNEL_NUMBER  => KERNEL_NUMBER,
        PADDING        => PADDING,
        STRIDE         => STRIDE
    )
    port map(
        clock        => clock,
        reset_n      => reset_n,
        i_sys_enable => i_sys_enable,
        i_data_valid => i_data_valid,
        i_data       => i_data,
        i_kernel     => i_kernel,
        i_bias       => i_bias,
        o_data       => o_data,
        o_data_valid => o_data_valid
    );

    i_bias <= (others => std_logic_vector(to_signed(-1, BITWIDTH)));

    -- Clock generation
    clock <= not clock after i_clk_period / 2;

    -------------------------------------------------------------------------------------
    -- TEST PROCESS
    -------------------------------------------------------------------------------------
    stimulus : process
        variable line_buffer : line;
    begin
        -- Reset the system
        reset_n      <= '0';
        i_data_valid <= '0';
        wait for i_clk_period;
        reset_n      <= '1';
        i_sys_enable <= '1';

        i_data(0) <= (
        (std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(62, 16))),
        (std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16))),
        (std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(66, 16))),
        (std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(251, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(60, 16))),
        (std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(60, 16))),
        (std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(254, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(59, 16))),
        (std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(16, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(253, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(12, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(251, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(31, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(22, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(12, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(24, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(65, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(60, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(62, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(65, 16))),
        (std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(28, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(68, 16))),
        (std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(12, 16)), std_logic_vector(to_signed(23, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(20, 16)), std_logic_vector(to_signed(16, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(70, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(26, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(32, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(26, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(31, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(19, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(16, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(56, 16))),
        (std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(19, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(13, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(251, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(29, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(62, 16))),
        (std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(21, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(19, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(68, 16))),
        (std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(69, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(252, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(70, 16))),
        (std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(31, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(254, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(71, 16))),
        (std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(62, 16))),
        (std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(253, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16))),
        (std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16))),
        (std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16))),
        (std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(72, 16))),
        (std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(75, 16))),
        (std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(72, 16))),
        (std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)))
        );
        i_data(1) <= (
        (std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(85, 16))),
        (std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(252, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16))),
        (std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(89, 16))),
        (std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(83, 16))),
        (std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(83, 16))),
        (std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(82, 16))),
        (std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(245, 16)), std_logic_vector(to_signed(254, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(16, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(252, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(13, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(13, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(251, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(32, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(23, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(254, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(12, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(254, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(24, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(28, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(88, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(83, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(85, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(90, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(88, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(249, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(31, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(31, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(25, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(32, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(93, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(20, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(30, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(84, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(13, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(12, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(79, 16))),
        (std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(85, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(91, 16))),
        (std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16))),
        (std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(85, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(85, 16))),
        (std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(88, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16))),
        (std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(252, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(89, 16))),
        (std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(87, 16))),
        (std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(82, 16))),
        (std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(77, 16))),
        (std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(224, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(226, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(72, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(238, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(75, 16))),
        (std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(72, 16))),
        (std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(231, 16)), std_logic_vector(to_signed(233, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(14, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16)))
        );
        i_data(2) <= (
        (std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16))),
        (std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(228, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(252, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16))),
        (std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(248, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(107, 16))),
        (std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(101, 16))),
        (std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(253, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(101, 16))),
        (std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(253, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(235, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(247, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(100, 16))),
        (std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(240, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(241, 16)), std_logic_vector(to_signed(255, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(232, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(20, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(229, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(19, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(239, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(217, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(244, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(230, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(237, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(223, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(24, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(107, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(222, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(22, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(29, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(106, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(101, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(108, 16))),
        (std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(242, 16)), std_logic_vector(to_signed(243, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(225, 16)), std_logic_vector(to_signed(250, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(106, 16))),
        (std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(234, 16)), std_logic_vector(to_signed(236, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(28, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(16, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(105, 16))),
        (std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(32, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16))),
        (std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(33, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(28, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(109, 16))),
        (std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(13, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(32, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(27, 16)), std_logic_vector(to_signed(221, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(22, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(111, 16))),
        (std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(251, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(28, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(18, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16))),
        (std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(246, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(25, 16)), std_logic_vector(to_signed(35, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(97, 16))),
        (std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(15, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(25, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(25, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(103, 16))),
        (std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16))),
        (std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(109, 16))),
        (std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(40, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(107, 16))),
        (std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(102, 16))),
        (std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(219, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(30, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(102, 16))),
        (std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(214, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(36, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(103, 16))),
        (std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(216, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(107, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(104, 16))),
        (std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(211, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(37, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(103, 16))),
        (std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(34, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(227, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16))),
        (std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(199, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(67, 16))),
        (std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(195, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(70, 16))),
        (std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(44, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(170, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(205, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(207, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(41, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(213, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(43, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(206, 16)), std_logic_vector(to_signed(215, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(188, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(76, 16))),
        (std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(174, 16)), std_logic_vector(to_signed(169, 16)), std_logic_vector(to_signed(171, 16)), std_logic_vector(to_signed(163, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(189, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(198, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(39, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(172, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(200, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(197, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(42, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(191, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(184, 16)), std_logic_vector(to_signed(194, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(48, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(209, 16)), std_logic_vector(to_signed(212, 16)), std_logic_vector(to_signed(196, 16)), std_logic_vector(to_signed(186, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(99, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(208, 16)), std_logic_vector(to_signed(203, 16)), std_logic_vector(to_signed(187, 16)), std_logic_vector(to_signed(179, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(193, 16)), std_logic_vector(to_signed(156, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(72, 16))),
        (std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(49, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(201, 16)), std_logic_vector(to_signed(210, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(3, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(10, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(164, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(166, 16)), std_logic_vector(to_signed(104, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(220, 16)), std_logic_vector(to_signed(180, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(12, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(17, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(45, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(190, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(204, 16)), std_logic_vector(to_signed(218, 16)), std_logic_vector(to_signed(176, 16)), std_logic_vector(to_signed(177, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(175, 16)), std_logic_vector(to_signed(185, 16)), std_logic_vector(to_signed(165, 16)), std_logic_vector(to_signed(181, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(102, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(202, 16)), std_logic_vector(to_signed(192, 16)), std_logic_vector(to_signed(182, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(173, 16)), std_logic_vector(to_signed(183, 16)), std_logic_vector(to_signed(178, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(167, 16)), std_logic_vector(to_signed(159, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(97, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(51, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(155, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(6, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(38, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(11, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(47, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(52, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(74, 16))),
        (std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(125, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(46, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(162, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(127, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(55, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(60, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(158, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(168, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(161, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(106, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(100, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(110, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(129, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(95, 16)), std_logic_vector(to_signed(92, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(152, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(126, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(160, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(76, 16)), std_logic_vector(to_signed(136, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(83, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(59, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(61, 16)), std_logic_vector(to_signed(65, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(121, 16)), std_logic_vector(to_signed(108, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(101, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(116, 16)), std_logic_vector(to_signed(150, 16)), std_logic_vector(to_signed(142, 16)), std_logic_vector(to_signed(135, 16)), std_logic_vector(to_signed(154, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(138, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(134, 16)), std_logic_vector(to_signed(131, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(149, 16)), std_logic_vector(to_signed(139, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(67, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(69, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(103, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(50, 16)), std_logic_vector(to_signed(79, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(93, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(62, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(96, 16)), std_logic_vector(to_signed(94, 16)), std_logic_vector(to_signed(73, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(109, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(118, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(124, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(140, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(153, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(133, 16)), std_logic_vector(to_signed(157, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(82, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(54, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(80, 16)), std_logic_vector(to_signed(70, 16)), std_logic_vector(to_signed(56, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16))),
        (std_logic_vector(to_signed(68, 16)), std_logic_vector(to_signed(53, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(58, 16)), std_logic_vector(to_signed(57, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(88, 16)), std_logic_vector(to_signed(75, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(81, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(63, 16)), std_logic_vector(to_signed(112, 16)), std_logic_vector(to_signed(117, 16)), std_logic_vector(to_signed(123, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(113, 16)), std_logic_vector(to_signed(119, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(115, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(122, 16)), std_logic_vector(to_signed(111, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(144, 16)), std_logic_vector(to_signed(137, 16)), std_logic_vector(to_signed(147, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(146, 16)), std_logic_vector(to_signed(148, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(151, 16)), std_logic_vector(to_signed(143, 16)), std_logic_vector(to_signed(145, 16)), std_logic_vector(to_signed(64, 16)), std_logic_vector(to_signed(72, 16)), std_logic_vector(to_signed(141, 16)), std_logic_vector(to_signed(114, 16)), std_logic_vector(to_signed(132, 16)), std_logic_vector(to_signed(130, 16)), std_logic_vector(to_signed(120, 16)), std_logic_vector(to_signed(105, 16)), std_logic_vector(to_signed(128, 16)), std_logic_vector(to_signed(74, 16)), std_logic_vector(to_signed(78, 16)), std_logic_vector(to_signed(77, 16)), std_logic_vector(to_signed(66, 16)), std_logic_vector(to_signed(98, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(89, 16)), std_logic_vector(to_signed(85, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(84, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(87, 16)), std_logic_vector(to_signed(90, 16)), std_logic_vector(to_signed(86, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(91, 16)), std_logic_vector(to_signed(71, 16)), std_logic_vector(to_signed(73, 16)))
        );

        -- FILTER EDGE
        i_kernel(0)(0) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)))
        );
        i_kernel(0)(1) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)))
        );
        i_kernel(0)(2) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(8, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)))
        );

        -- FILTER EMBOSS
        i_kernel(1)(0) <= (
        (std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(2, 16)))
        );
        i_kernel(1)(1) <= (
        (std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(2, 16)))
        );
        i_kernel(1)(2) <= (
        (std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(2, 16)))
        );

        -- FILTER IDENTITY
        i_kernel(2)(0) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)))
        );
        i_kernel(2)(1) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)))
        );
        i_kernel(2)(2) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)))
        );

        -- FILTER LAPLACIAN DIAG
        i_kernel(3)(0) <= (
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(-8, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(3)(1) <= (
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(-8, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(3)(2) <= (
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(-8, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)))
        );

        -- FILTER PREWITT X AXIS
        i_kernel(4)(0) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(4)(1) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(4)(2) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)))
        );

        -- FILTER PREWITT Y AXIS
        i_kernel(5)(0) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(5)(1) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(5)(2) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(1, 16)))
        );

        -- FILTER RANDOM
        i_kernel(6)(0) <= (
        (std_logic_vector(to_signed(-10, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(-9, 16))),
        (std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(-7, 16))),
        (std_logic_vector(to_signed(-4, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(-4, 16)))
        );
        i_kernel(6)(1) <= (
        (std_logic_vector(to_signed(-10, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(-9, 16))),
        (std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(-7, 16))),
        (std_logic_vector(to_signed(-4, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(-4, 16)))
        );
        i_kernel(6)(2) <= (
        (std_logic_vector(to_signed(-10, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(-9, 16))),
        (std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(7, 16)), std_logic_vector(to_signed(-7, 16))),
        (std_logic_vector(to_signed(-4, 16)), std_logic_vector(to_signed(9, 16)), std_logic_vector(to_signed(-4, 16)))
        );

        -- FILTER RIDGE
        i_kernel(7)(0) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)))
        );
        i_kernel(7)(1) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)))
        );
        i_kernel(7)(2) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(4, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)))
        );

        -- FILTER SHARP
        i_kernel(8)(0) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)))
        );
        i_kernel(8)(1) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)))
        );
        i_kernel(8)(2) <= (
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(5, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)))
        );

        -- FILTER SOBEL X
        i_kernel(9)(0) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(2, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(9)(1) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(2, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(9)(2) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16))),
        (std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(2, 16))),
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(1, 16)))
        );

        -- FILTER SOBEL Y
        i_kernel(10)(0) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(10)(1) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(1, 16)))
        );
        i_kernel(10)(2) <= (
        (std_logic_vector(to_signed(-1, 16)), std_logic_vector(to_signed(-2, 16)), std_logic_vector(to_signed(-1, 16))),
        (std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16)), std_logic_vector(to_signed(0, 16))),
        (std_logic_vector(to_signed(1, 16)), std_logic_vector(to_signed(2, 16)), std_logic_vector(to_signed(1, 16)))
        );

        -- FILTER BLUR * 1000
        i_kernel(11)(0) <= (
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16))),
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16))),
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)))
        );
        i_kernel(11)(1) <= (
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16))),
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16))),
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)))
        );
        i_kernel(11)(2) <= (
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16))),
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16))),
        (std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)), std_logic_vector(to_signed(1111, 16)))
        );

        -- GAUSSIAN FITLER * 1000
        i_kernel(12)(0) <= (
        (std_logic_vector(to_signed(625, 16)), std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(625, 16))),
        (std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(2500, 16)), std_logic_vector(to_signed(1250, 16))),
        (std_logic_vector(to_signed(625, 16)), std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(625, 16)))
        );
        i_kernel(12)(1) <= (
        (std_logic_vector(to_signed(625, 16)), std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(625, 16))),
        (std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(2500, 16)), std_logic_vector(to_signed(1250, 16))),
        (std_logic_vector(to_signed(625, 16)), std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(625, 16)))
        );
        i_kernel(12)(2) <= (
        (std_logic_vector(to_signed(625, 16)), std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(625, 16))),
        (std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(2500, 16)), std_logic_vector(to_signed(1250, 16))),
        (std_logic_vector(to_signed(625, 16)), std_logic_vector(to_signed(1250, 16)), std_logic_vector(to_signed(625, 16)))
        );

        wait for i_clk_period/2;
        i_data_valid <= '1';
        wait for i_clk_period;
        i_data_valid <= '0';

        -- Open the file
        file_open(output_file, "conv2d_output_results.txt", write_mode);

        -- Wait for output to be valid and write to file
        wait until o_data_valid = '1';
        for k in 0 to KERNEL_NUMBER - 1 loop
            for i in ((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1) downto 0 loop
                for j in ((INPUT_SIZE + 2 * PADDING - KERNEL_SIZE)/STRIDE + 1 - 1) downto 0 loop
                    write(line_buffer, o_data(k)(i)(j));
                    writeline(output_file, line_buffer);
                end loop;
            end loop;
        end loop;

        -- Close the file
        file_close(output_file);

        -- End simulation
        wait;

    end process stimulus;
end conv2d_tb_arch;

configuration conv2d_tb_conf of conv2d_tb is
    for conv2d_tb_arch
        for UUT : conv2d
            use configuration LIB_RTL.conv2d_fc_conf;
        end for;
    end for;
end configuration conv2d_tb_conf;